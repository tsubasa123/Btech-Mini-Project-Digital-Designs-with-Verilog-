module VGA_Control (clock, reset, ::);
